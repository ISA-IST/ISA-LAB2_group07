	SIGNAL sum_0, c_out_0: STD_LOGIC_VECTOR (51 downto 0);
	SIGNAL sum_1, c_out_1: STD_LOGIC_VECTOR (115 downto 0);
	SIGNAL sum_2, c_out_2: STD_LOGIC_VECTOR (128 downto 0);
	SIGNAL sum_3, c_out_3: STD_LOGIC_VECTOR (105 downto 0);
	SIGNAL sum_4, c_out_4: STD_LOGIC_VECTOR (58 downto 0);
	SIGNAL sum_5, c_out_5: STD_LOGIC_VECTOR (61 downto 0);
	SIGNAL sum_6, c_out_6: STD_LOGIC;

BEGIN

