
	HA_6 : HA port map (A=>pp0(0), B=>s(0), S=>sum_6, C_out=>c_out_6);

	addend1_out <= sum_5(61) & sum_5(60) & sum_5(59) & sum_5(58) & sum_5(57) & sum_5(56) & sum_5(55) & sum_5(54) & sum_5(53) & sum_5(52) & sum_5(51) & sum_5(50) & sum_5(49) & sum_5(48) & sum_5(47) & sum_5(46) & sum_5(45) & sum_5(44) & sum_5(43) & sum_5(42) & sum_5(41) & sum_5(40) & sum_5(39) & sum_5(38) & sum_5(37) & sum_5(36) & sum_5(35) & sum_5(34) & sum_5(33) & sum_5(32) & sum_5(31) & sum_5(30) & sum_5(29) & sum_5(28) & sum_5(27) & sum_5(26) & sum_5(25) & sum_5(24) & sum_5(23) & sum_5(22) & sum_5(21) & sum_5(20) & sum_5(19) & sum_5(18) & sum_5(17) & sum_5(16) & sum_5(15) & sum_5(14) & sum_5(13) & sum_5(12) & sum_5(11) & sum_5(10) & sum_5(9) & sum_5(8) & sum_5(7) & sum_5(6) & sum_5(5) & sum_5(4) & sum_5(3) & sum_5(2) & sum_5(1) & sum_5(0) & c_out_6;

	addend2_out <= c_out_5(60) & c_out_5(59) & c_out_5(58) & c_out_5(57) & c_out_5(56) & c_out_5(55) & c_out_5(54) & c_out_5(53) & c_out_5(52) & c_out_5(51) & c_out_5(50) & c_out_5(49) & c_out_5(48) & c_out_5(47) & c_out_5(46) & c_out_5(45) & c_out_5(44) & c_out_5(43) & c_out_5(42) & c_out_5(41) & c_out_5(40) & c_out_5(39) & c_out_5(38) & c_out_5(37) & c_out_5(36) & c_out_5(35) & c_out_5(34) & c_out_5(33) & c_out_5(32) & c_out_5(31) & c_out_5(30) & c_out_5(29) & c_out_5(28) & c_out_5(27) & c_out_5(26) & c_out_5(25) & c_out_5(24) & c_out_5(23) & c_out_5(22) & c_out_5(21) & c_out_5(20) & c_out_5(19) & c_out_5(18) & c_out_5(17) & c_out_5(16) & c_out_5(15) & c_out_5(14) & c_out_5(13) & c_out_5(12) & c_out_5(11) & c_out_5(10) & c_out_5(9) & c_out_5(8) & c_out_5(7) & c_out_5(6) & c_out_5(5) & c_out_5(4) & c_out_5(3) & c_out_5(2) & c_out_5(1) & c_out_5(0) & pp0(2) & pp0(1);

	M_lsb <= sum_6;

END struct;