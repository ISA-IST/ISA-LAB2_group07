	SIGNAL : sum_0, c_out_0: std_logic_vector (51 downto 0);
	SIGNAL : sum_1, c_out_1: std_logic_vector (115 downto 0);
	SIGNAL : sum_2, c_out_2: std_logic_vector (128 downto 0);
	SIGNAL : sum_3, c_out_3: std_logic_vector (105 downto 0);
	SIGNAL : sum_4, c_out_4: std_logic_vector (58 downto 0);
	SIGNAL : sum_5, c_out_5: std_logic_vector (61 downto 0);
	SIGNAL : sum_6, c_out_6;

BEGIN

