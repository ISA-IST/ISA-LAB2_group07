library verilog;
use verilog.vl_types.all;
entity tb_mult_pipe is
end tb_mult_pipe;
