library verilog;
use verilog.vl_types.all;
entity tb_MBE_mult is
end tb_MBE_mult;
